library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

-- Entity declaration for the alarm clock
entity AlarmClock is
    Port (
        clk         : in STD_LOGIC;     -- Input clock (e.g., 50 MHz)
        reset       : in STD_LOGIC;     -- Asynchronous reset
        set_alarm   : in STD_LOGIC;     -- Set alarm signal
        set_time    : in STD_LOGIC;     -- Set time signal
        alarm_time  : in STD_LOGIC_VECTOR(7 downto 0); -- Alarm time (hour, minute)
        current_time: out STD_LOGIC_VECTOR(7 downto 0); -- Current time (hour, minute)
        alarm       : out STD_LOGIC      -- Alarm output
    );
end AlarmClock;

-- Architecture definition for the alarm clock
architecture Behavioral of AlarmClock is
    signal clk_div  : STD_LOGIC := '0';  -- Divided clock signal (1 Hz pulse)
    signal sec_count: integer := 0;      -- Second counter
    signal min_count: integer := 0;      -- Minute counter
    signal hr_count : integer := 0;      -- Hour counter
    signal alarm_time_reg : STD_LOGIC_VECTOR(7 downto 0) := (others => '0');
    signal alarm_match : STD_LOGIC := '0';

    -- Clock division process
    process(clk, reset)
    begin
        if reset = '1' then
            clk_div <= '0';
            sec_count <= 0;
        elsif rising_edge(clk) then
            if sec_count = 49999999 then  -- Assuming clk is 50 MHz
                clk_div <= not clk_div;
                sec_count <= 0;
            else
                sec_count <= sec_count + 1;
            end if;
        end if;
    end process;

    -- Time counter process
    process(clk_div, reset)
    begin
        if reset = '1' then
            min_count <= 0;
            hr_count <= 0;
        elsif rising_edge(clk_div) then
            if min_count = 59 then
                min_count <= 0;
                if hr_count = 23 then
                    hr_count <= 0;
                else
                    hr_count <= hr_count + 1;
                end if;
            else
                min_count <= min_count + 1;
            end if;
        end if;
    end process;

    -- Alarm comparison process
    process(set_alarm, clk_div, reset)
    begin
        if reset = '1' then
            alarm_time_reg <= (others => '0');
            alarm_match <= '0';
        elsif set_alarm = '1' then
            alarm_time_reg <= alarm_time;
        else
            if (std_logic_vector(to_unsigned(hr_count, 4)) & std_logic_vector(to_unsigned(min_count, 4))) = alarm_time_reg then
                alarm_match <= '1';
            else
                alarm_match <= '0';
            end if;
        end if;
    end process;

    -- Output assignment
    current_time <= std_logic_vector(to_unsigned(hr_count, 4)) & std_logic_vector(to_unsigned(min_count, 4));
    alarm <= alarm_match;

end Behavioral;













































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































--Akhil Rai
